/*************************************************************************
   > File Name:     defines.svh
   > Description:   This File contains the macro definitions.
   > Author:        Noman Rafiq
   > Modified:      Dec 10, 2024
   > Mail:          noman.rafiq@10xengineers.ai
   ---------------------------------------------------------------
   Copyright   (c)2024 10xEngineers
   ---------------------------------------------------------------
************************************************************************/  

  // Source and Destination Addresses for Read/Writes
  `define SRC_ADDR 32'h0;
  `define DST_ADDR 32'h0;