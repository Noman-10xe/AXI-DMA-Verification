// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
`ifndef MEM_MODEL_PKG
`define MEM_MODEL_PKG

package mem_model_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "dv_macros.svh"
  `include "mem_model.sv"

endpackage
`endif